module led(
    input wire sclk

);

endmodule